-- nios.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios is
	port (
		amwr_address      : in    std_logic_vector(31 downto 0) := (others => '0'); --     amwr.address
		amwr_byteenable   : in    std_logic_vector(3 downto 0)  := (others => '0'); --         .byteenable
		amwr_write        : in    std_logic                     := '0';             --         .write
		amwr_writedata    : in    std_logic_vector(31 downto 0) := (others => '0'); --         .writedata
		amwr_waitrequest  : out   std_logic;                                        --         .waitrequest
		amwr_burstcount   : in    std_logic_vector(7 downto 0)  := (others => '0'); --         .burstcount
		as_pdm_address    : out   std_logic_vector(9 downto 0);                     --   as_pdm.address
		as_pdm_read       : out   std_logic;                                        --         .read
		as_pdm_readdata   : in    std_logic_vector(31 downto 0) := (others => '0'); --         .readdata
		as_pdm_write      : out   std_logic;                                        --         .write
		as_pdm_writedata  : out   std_logic_vector(31 downto 0);                    --         .writedata
		as_pdm_byteenable : out   std_logic_vector(3 downto 0);                     --         .byteenable
		as_pdm_chipselect : out   std_logic;                                        --         .chipselect
		button_export     : in    std_logic_vector(3 downto 0)  := (others => '0'); --   button.export
		clk_clk           : in    std_logic                     := '0';             --      clk.clk
		deb_export        : out   std_logic_vector(7 downto 0);                     --      deb.export
		ftdi_rdn          : out   std_logic;                                        --     ftdi.rdn
		ftdi_resetn       : out   std_logic;                                        --         .resetn
		ftdi_rxdata       : in    std_logic_vector(7 downto 0)  := (others => '0'); --         .rxdata
		ftdi_rxfn         : in    std_logic                     := '0';             --         .rxfn
		ftdi_txdata       : out   std_logic_vector(7 downto 0);                     --         .txdata
		ftdi_txdata_oe    : out   std_logic;                                        --         .txdata_oe
		ftdi_txen         : in    std_logic                     := '0';             --         .txen
		ftdi_wr           : out   std_logic;                                        --         .wr
		lcd_cs            : out   std_logic;                                        --      lcd.cs
		lcd_dc            : out   std_logic;                                        --         .dc
		lcd_rstn          : out   std_logic;                                        --         .rstn
		lcd_sclk          : out   std_logic;                                        --         .sclk
		lcd_sdata         : out   std_logic;                                        --         .sdata
		led_export        : out   std_logic_vector(7 downto 0);                     --      led.export
		log_clk           : out   std_logic;                                        --      log.clk
		pdm_clk           : out   std_logic;                                        --      pdm.clk
		pll_lock_export   : out   std_logic;                                        -- pll_lock.export
		reset_reset_n     : in    std_logic                     := '0';             --    reset.reset_n
		sd_clk            : out   std_logic;                                        --       sd.clk
		sdram_addr        : out   std_logic_vector(11 downto 0);                    --    sdram.addr
		sdram_ba          : out   std_logic_vector(1 downto 0);                     --         .ba
		sdram_cas_n       : out   std_logic;                                        --         .cas_n
		sdram_cke         : out   std_logic;                                        --         .cke
		sdram_cs_n        : out   std_logic;                                        --         .cs_n
		sdram_dq          : inout std_logic_vector(15 downto 0) := (others => '0'); --         .dq
		sdram_dqm         : out   std_logic_vector(1 downto 0);                     --         .dqm
		sdram_ras_n       : out   std_logic;                                        --         .ras_n
		sdram_we_n        : out   std_logic;                                        --         .we_n
		sflash_dclk       : out   std_logic;                                        --   sflash.dclk
		sflash_sce        : out   std_logic;                                        --         .sce
		sflash_sdo        : out   std_logic;                                        --         .sdo
		sflash_data0      : in    std_logic                     := '0';             --         .data0
		sys_clk           : out   std_logic                                         --      sys.clk
	);
end entity nios;

architecture rtl of nios is
	component nios_DEBport is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios_DEBport;

	component ili9341_spi16 is
		port (
			clk     : in  std_logic                     := 'X';             -- clk
			reset_n : in  std_logic                     := 'X';             -- reset_n
			address : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			ben     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			sel     : in  std_logic                     := 'X';             -- chipselect
			wr      : in  std_logic                     := 'X';             -- write
			wrdata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			waitreq : out std_logic;                                        -- waitrequest
			cs      : out std_logic;                                        -- cs
			dc      : out std_logic;                                        -- dc
			rstn    : out std_logic;                                        -- rstn
			sclk    : out std_logic;                                        -- sclk
			sdata   : out std_logic                                         -- sdata
		);
	end component ili9341_spi16;

	component nios_button is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component nios_button;

	component nios_dma is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			system_reset_n     : in  std_logic                     := 'X';             -- reset_n
			dma_ctl_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			dma_ctl_chipselect : in  std_logic                     := 'X';             -- chipselect
			dma_ctl_readdata   : out std_logic_vector(23 downto 0);                    -- readdata
			dma_ctl_write_n    : in  std_logic                     := 'X';             -- write_n
			dma_ctl_writedata  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- writedata
			dma_ctl_irq        : out std_logic;                                        -- irq
			read_address       : out std_logic_vector(23 downto 0);                    -- address
			read_chipselect    : out std_logic;                                        -- chipselect
			read_read_n        : out std_logic;                                        -- read_n
			read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			write_address      : out std_logic_vector(23 downto 0);                    -- address
			write_chipselect   : out std_logic;                                        -- chipselect
			write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			write_write_n      : out std_logic;                                        -- write_n
			write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			write_byteenable   : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component nios_dma;

	component nios_dma_LCD is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			system_reset_n     : in  std_logic                     := 'X';             -- reset_n
			dma_ctl_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			dma_ctl_chipselect : in  std_logic                     := 'X';             -- chipselect
			dma_ctl_readdata   : out std_logic_vector(23 downto 0);                    -- readdata
			dma_ctl_write_n    : in  std_logic                     := 'X';             -- write_n
			dma_ctl_writedata  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- writedata
			dma_ctl_irq        : out std_logic;                                        -- irq
			read_address       : out std_logic_vector(23 downto 0);                    -- address
			read_chipselect    : out std_logic;                                        -- chipselect
			read_read_n        : out std_logic;                                        -- read_n
			read_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			write_address      : out std_logic_vector(23 downto 0);                    -- address
			write_chipselect   : out std_logic;                                        -- chipselect
			write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			write_write_n      : out std_logic;                                        -- write_n
			write_writedata    : out std_logic_vector(15 downto 0);                    -- writedata
			write_byteenable   : out std_logic_vector(1 downto 0)                      -- byteenable
		);
	end component nios_dma_LCD;

	component ft245if2 is
		port (
			address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			ben          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			rd           : in  std_logic                     := 'X';             -- read
			rddata       : out std_logic_vector(31 downto 0);                    -- readdata
			sel          : in  std_logic                     := 'X';             -- chipselect
			waitreq      : out std_logic;                                        -- waitrequest
			wr           : in  std_logic                     := 'X';             -- write
			wrdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clk          : in  std_logic                     := 'X';             -- clk
			ft_rdn       : out std_logic;                                        -- rdn
			ft_resetn    : out std_logic;                                        -- resetn
			ft_rxdata    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rxdata
			ft_rxfn      : in  std_logic                     := 'X';             -- rxfn
			ft_txdata    : out std_logic_vector(7 downto 0);                     -- txdata
			ft_txdata_oe : out std_logic;                                        -- txdata_oe
			ft_txen      : in  std_logic                     := 'X';             -- txen
			ft_wr        : out std_logic;                                        -- wr
			irq          : out std_logic;                                        -- irq
			reset_n      : in  std_logic                     := 'X'              -- reset_n
		);
	end component ft245if2;

	component nios_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_jtag_uart;

	component nios_nios2_gen2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(23 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(23 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_nios2_gen2;

	component altera_onchip_flash is
		generic (
			INIT_FILENAME                       : string  := "";
			INIT_FILENAME_SIM                   : string  := "";
			DEVICE_FAMILY                       : string  := "Unknown";
			PART_NAME                           : string  := "Unknown";
			DEVICE_ID                           : string  := "Unknown";
			SECTOR1_START_ADDR                  : integer := 0;
			SECTOR1_END_ADDR                    : integer := 0;
			SECTOR2_START_ADDR                  : integer := 0;
			SECTOR2_END_ADDR                    : integer := 0;
			SECTOR3_START_ADDR                  : integer := 0;
			SECTOR3_END_ADDR                    : integer := 0;
			SECTOR4_START_ADDR                  : integer := 0;
			SECTOR4_END_ADDR                    : integer := 0;
			SECTOR5_START_ADDR                  : integer := 0;
			SECTOR5_END_ADDR                    : integer := 0;
			MIN_VALID_ADDR                      : integer := 0;
			MAX_VALID_ADDR                      : integer := 0;
			MIN_UFM_VALID_ADDR                  : integer := 0;
			MAX_UFM_VALID_ADDR                  : integer := 0;
			SECTOR1_MAP                         : integer := 0;
			SECTOR2_MAP                         : integer := 0;
			SECTOR3_MAP                         : integer := 0;
			SECTOR4_MAP                         : integer := 0;
			SECTOR5_MAP                         : integer := 0;
			ADDR_RANGE1_END_ADDR                : integer := 0;
			ADDR_RANGE2_END_ADDR                : integer := 0;
			ADDR_RANGE1_OFFSET                  : integer := 0;
			ADDR_RANGE2_OFFSET                  : integer := 0;
			ADDR_RANGE3_OFFSET                  : integer := 0;
			AVMM_DATA_ADDR_WIDTH                : integer := 19;
			AVMM_DATA_DATA_WIDTH                : integer := 32;
			AVMM_DATA_BURSTCOUNT_WIDTH          : integer := 4;
			SECTOR_READ_PROTECTION_MODE         : integer := 31;
			FLASH_SEQ_READ_DATA_COUNT           : integer := 2;
			FLASH_ADDR_ALIGNMENT_BITS           : integer := 1;
			FLASH_READ_CYCLE_MAX_INDEX          : integer := 4;
			FLASH_RESET_CYCLE_MAX_INDEX         : integer := 29;
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  : integer := 112;
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX : integer := 40603248;
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX : integer := 35382;
			PARALLEL_MODE                       : boolean := true;
			READ_AND_WRITE_MODE                 : boolean := true;
			WRAPPING_BURST_MODE                 : boolean := false;
			IS_DUAL_BOOT                        : string  := "False";
			IS_ERAM_SKIP                        : string  := "False";
			IS_COMPRESSED_IMAGE                 : string  := "False"
		);
		port (
			clock                   : in  std_logic                     := 'X';             -- clk
			reset_n                 : in  std_logic                     := 'X';             -- reset_n
			avmm_data_addr          : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			avmm_data_read          : in  std_logic                     := 'X';             -- read
			avmm_data_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_data_write         : in  std_logic                     := 'X';             -- write
			avmm_data_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avmm_data_waitrequest   : out std_logic;                                        -- waitrequest
			avmm_data_readdatavalid : out std_logic;                                        -- readdatavalid
			avmm_data_burstcount    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			avmm_csr_addr           : in  std_logic                     := 'X';             -- address
			avmm_csr_read           : in  std_logic                     := 'X';             -- read
			avmm_csr_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_csr_write          : in  std_logic                     := 'X';             -- write
			avmm_csr_readdata       : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component altera_onchip_flash;

	component nios_pll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component nios_pll;

	component nios_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component nios_sdram;

	component nios_serialflash is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read_n     : in  std_logic                     := 'X';             -- read_n
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			irq        : out std_logic;                                        -- irq
			dclk       : out std_logic;                                        -- export
			sce        : out std_logic;                                        -- export
			sdo        : out std_logic;                                        -- export
			data0      : in  std_logic                     := 'X'              -- export
		);
	end component nios_serialflash;

	component nios_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_sys_clk_timer;

	component nios_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios_sysid;

	component nios_mm_interconnect_0 is
		port (
			pll_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			av_wr_master_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_uart_reset_reset_bridge_in_reset_reset           : in  std_logic                     := 'X';             -- reset
			nios2_gen2_reset_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			av_wr_master_0_avalon_master_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_wr_master_0_avalon_master_waitrequest              : out std_logic;                                        -- waitrequest
			av_wr_master_0_avalon_master_burstcount               : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			av_wr_master_0_avalon_master_byteenable               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_wr_master_0_avalon_master_write                    : in  std_logic                     := 'X';             -- write
			av_wr_master_0_avalon_master_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dma_read_master_address                               : in  std_logic_vector(23 downto 0) := (others => 'X'); -- address
			dma_read_master_waitrequest                           : out std_logic;                                        -- waitrequest
			dma_read_master_chipselect                            : in  std_logic                     := 'X';             -- chipselect
			dma_read_master_read                                  : in  std_logic                     := 'X';             -- read
			dma_read_master_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			dma_read_master_readdatavalid                         : out std_logic;                                        -- readdatavalid
			dma_write_master_address                              : in  std_logic_vector(23 downto 0) := (others => 'X'); -- address
			dma_write_master_waitrequest                          : out std_logic;                                        -- waitrequest
			dma_write_master_byteenable                           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			dma_write_master_chipselect                           : in  std_logic                     := 'X';             -- chipselect
			dma_write_master_write                                : in  std_logic                     := 'X';             -- write
			dma_write_master_writedata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dma_LCD_read_master_address                           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- address
			dma_LCD_read_master_waitrequest                       : out std_logic;                                        -- waitrequest
			dma_LCD_read_master_chipselect                        : in  std_logic                     := 'X';             -- chipselect
			dma_LCD_read_master_read                              : in  std_logic                     := 'X';             -- read
			dma_LCD_read_master_readdata                          : out std_logic_vector(15 downto 0);                    -- readdata
			dma_LCD_read_master_readdatavalid                     : out std_logic;                                        -- readdatavalid
			dma_LCD_write_master_address                          : in  std_logic_vector(23 downto 0) := (others => 'X'); -- address
			dma_LCD_write_master_waitrequest                      : out std_logic;                                        -- waitrequest
			dma_LCD_write_master_byteenable                       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			dma_LCD_write_master_chipselect                       : in  std_logic                     := 'X';             -- chipselect
			dma_LCD_write_master_write                            : in  std_logic                     := 'X';             -- write
			dma_LCD_write_master_writedata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_data_master_address                        : in  std_logic_vector(23 downto 0) := (others => 'X'); -- address
			nios2_gen2_data_master_waitrequest                    : out std_logic;                                        -- waitrequest
			nios2_gen2_data_master_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_data_master_read                           : in  std_logic                     := 'X';             -- read
			nios2_gen2_data_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_data_master_write                          : in  std_logic                     := 'X';             -- write
			nios2_gen2_data_master_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_data_master_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_instruction_master_address                 : in  std_logic_vector(23 downto 0) := (others => 'X'); -- address
			nios2_gen2_instruction_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_gen2_instruction_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_gen2_instruction_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			button_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			button_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DEBport_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			DEBport_s1_write                                      : out std_logic;                                        -- write
			DEBport_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DEBport_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			DEBport_s1_chipselect                                 : out std_logic;                                        -- chipselect
			dma_control_port_slave_address                        : out std_logic_vector(2 downto 0);                     -- address
			dma_control_port_slave_write                          : out std_logic;                                        -- write
			dma_control_port_slave_readdata                       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- readdata
			dma_control_port_slave_writedata                      : out std_logic_vector(23 downto 0);                    -- writedata
			dma_control_port_slave_chipselect                     : out std_logic;                                        -- chipselect
			dma_LCD_control_port_slave_address                    : out std_logic_vector(2 downto 0);                     -- address
			dma_LCD_control_port_slave_write                      : out std_logic;                                        -- write
			dma_LCD_control_port_slave_readdata                   : in  std_logic_vector(23 downto 0) := (others => 'X'); -- readdata
			dma_LCD_control_port_slave_writedata                  : out std_logic_vector(23 downto 0);                    -- writedata
			dma_LCD_control_port_slave_chipselect                 : out std_logic;                                        -- chipselect
			ft245_avalon_slave_address                            : out std_logic_vector(2 downto 0);                     -- address
			ft245_avalon_slave_write                              : out std_logic;                                        -- write
			ft245_avalon_slave_read                               : out std_logic;                                        -- read
			ft245_avalon_slave_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ft245_avalon_slave_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			ft245_avalon_slave_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			ft245_avalon_slave_waitrequest                        : in  std_logic                     := 'X';             -- waitrequest
			ft245_avalon_slave_chipselect                         : out std_logic;                                        -- chipselect
			ILI9341SPI_a_slave_address                            : out std_logic_vector(1 downto 0);                     -- address
			ILI9341SPI_a_slave_write                              : out std_logic;                                        -- write
			ILI9341SPI_a_slave_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			ILI9341SPI_a_slave_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			ILI9341SPI_a_slave_waitrequest                        : in  std_logic                     := 'X';             -- waitrequest
			ILI9341SPI_a_slave_chipselect                         : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                     : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                      : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                : out std_logic;                                        -- chipselect
			LED_s1_address                                        : out std_logic_vector(1 downto 0);                     -- address
			LED_s1_write                                          : out std_logic;                                        -- write
			LED_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LED_s1_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			LED_s1_chipselect                                     : out std_logic;                                        -- chipselect
			nios2_gen2_debug_mem_slave_address                    : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_debug_mem_slave_write                      : out std_logic;                                        -- write
			nios2_gen2_debug_mem_slave_read                       : out std_logic;                                        -- read
			nios2_gen2_debug_mem_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_debug_mem_slave_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_debug_mem_slave_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_debug_mem_slave_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_debug_mem_slave_debugaccess                : out std_logic;                                        -- debugaccess
			onchip_flash_data_address                             : out std_logic_vector(12 downto 0);                    -- address
			onchip_flash_data_write                               : out std_logic;                                        -- write
			onchip_flash_data_read                                : out std_logic;                                        -- read
			onchip_flash_data_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_data_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_data_burstcount                          : out std_logic_vector(3 downto 0);                     -- burstcount
			onchip_flash_data_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			onchip_flash_data_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			pdm_s0_address                                        : out std_logic_vector(9 downto 0);                     -- address
			pdm_s0_write                                          : out std_logic;                                        -- write
			pdm_s0_read                                           : out std_logic;                                        -- read
			pdm_s0_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pdm_s0_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			pdm_s0_byteenable                                     : out std_logic_vector(3 downto 0);                     -- byteenable
			pdm_s0_chipselect                                     : out std_logic;                                        -- chipselect
			sdram_s1_address                                      : out std_logic_vector(21 downto 0);                    -- address
			sdram_s1_write                                        : out std_logic;                                        -- write
			sdram_s1_read                                         : out std_logic;                                        -- read
			sdram_s1_readdata                                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                    : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                                   : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                   : out std_logic;                                        -- chipselect
			serialflash_epcs_control_port_address                 : out std_logic_vector(8 downto 0);                     -- address
			serialflash_epcs_control_port_write                   : out std_logic;                                        -- write
			serialflash_epcs_control_port_read                    : out std_logic;                                        -- read
			serialflash_epcs_control_port_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			serialflash_epcs_control_port_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			serialflash_epcs_control_port_chipselect              : out std_logic;                                        -- chipselect
			sys_clk_timer_s1_address                              : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                                : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata                             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata                            : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect                           : out std_logic;                                        -- chipselect
			sysid_control_slave_address                           : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component nios_mm_interconnect_0;

	component nios_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_irq_mapper;

	component nios_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_rst_controller;

	component nios_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_rst_controller_001;

	signal pll_c0_clk                                                      : std_logic;                     -- pll:c0 -> [DEBport:clk, ILI9341SPI:clk, LED:clk, button:clk, dma:clk, dma_LCD:clk, ft245:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:pll_c0_clk, nios2_gen2:clk, onchip_flash:clock, rst_controller:clk, rst_controller_001:clk, sdram:clk, serialflash:clk, sys_clk_timer:clk, sysid:clock]
	signal nios2_gen2_debug_reset_request_reset                            : std_logic;                     -- nios2_gen2:debug_reset_request -> [mm_interconnect_0:av_wr_master_0_reset_sink_reset_bridge_in_reset_reset, nios2_gen2_debug_reset_request_reset:in, rst_controller:reset_in1]
	signal nios2_gen2_data_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	signal nios2_gen2_data_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	signal nios2_gen2_data_master_debugaccess                              : std_logic;                     -- nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	signal nios2_gen2_data_master_address                                  : std_logic_vector(23 downto 0); -- nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	signal nios2_gen2_data_master_byteenable                               : std_logic_vector(3 downto 0);  -- nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	signal nios2_gen2_data_master_read                                     : std_logic;                     -- nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	signal nios2_gen2_data_master_write                                    : std_logic;                     -- nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	signal nios2_gen2_data_master_writedata                                : std_logic_vector(31 downto 0); -- nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	signal nios2_gen2_instruction_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	signal nios2_gen2_instruction_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	signal nios2_gen2_instruction_master_address                           : std_logic_vector(23 downto 0); -- nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	signal nios2_gen2_instruction_master_read                              : std_logic;                     -- nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	signal dma_read_master_chipselect                                      : std_logic;                     -- dma:read_chipselect -> mm_interconnect_0:dma_read_master_chipselect
	signal dma_read_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:dma_read_master_readdata -> dma:read_readdata
	signal dma_read_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:dma_read_master_waitrequest -> dma:read_waitrequest
	signal dma_read_master_address                                         : std_logic_vector(23 downto 0); -- dma:read_address -> mm_interconnect_0:dma_read_master_address
	signal dma_read_master_read                                            : std_logic;                     -- dma:read_read_n -> dma_read_master_read:in
	signal dma_read_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:dma_read_master_readdatavalid -> dma:read_readdatavalid
	signal dma_lcd_read_master_chipselect                                  : std_logic;                     -- dma_LCD:read_chipselect -> mm_interconnect_0:dma_LCD_read_master_chipselect
	signal dma_lcd_read_master_readdata                                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:dma_LCD_read_master_readdata -> dma_LCD:read_readdata
	signal dma_lcd_read_master_waitrequest                                 : std_logic;                     -- mm_interconnect_0:dma_LCD_read_master_waitrequest -> dma_LCD:read_waitrequest
	signal dma_lcd_read_master_address                                     : std_logic_vector(23 downto 0); -- dma_LCD:read_address -> mm_interconnect_0:dma_LCD_read_master_address
	signal dma_lcd_read_master_read                                        : std_logic;                     -- dma_LCD:read_read_n -> dma_lcd_read_master_read:in
	signal dma_lcd_read_master_readdatavalid                               : std_logic;                     -- mm_interconnect_0:dma_LCD_read_master_readdatavalid -> dma_LCD:read_readdatavalid
	signal dma_write_master_chipselect                                     : std_logic;                     -- dma:write_chipselect -> mm_interconnect_0:dma_write_master_chipselect
	signal dma_write_master_waitrequest                                    : std_logic;                     -- mm_interconnect_0:dma_write_master_waitrequest -> dma:write_waitrequest
	signal dma_write_master_address                                        : std_logic_vector(23 downto 0); -- dma:write_address -> mm_interconnect_0:dma_write_master_address
	signal dma_write_master_byteenable                                     : std_logic_vector(3 downto 0);  -- dma:write_byteenable -> mm_interconnect_0:dma_write_master_byteenable
	signal dma_write_master_write                                          : std_logic;                     -- dma:write_write_n -> dma_write_master_write:in
	signal dma_write_master_writedata                                      : std_logic_vector(31 downto 0); -- dma:write_writedata -> mm_interconnect_0:dma_write_master_writedata
	signal dma_lcd_write_master_chipselect                                 : std_logic;                     -- dma_LCD:write_chipselect -> mm_interconnect_0:dma_LCD_write_master_chipselect
	signal dma_lcd_write_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:dma_LCD_write_master_waitrequest -> dma_LCD:write_waitrequest
	signal dma_lcd_write_master_address                                    : std_logic_vector(23 downto 0); -- dma_LCD:write_address -> mm_interconnect_0:dma_LCD_write_master_address
	signal dma_lcd_write_master_byteenable                                 : std_logic_vector(1 downto 0);  -- dma_LCD:write_byteenable -> mm_interconnect_0:dma_LCD_write_master_byteenable
	signal dma_lcd_write_master_write                                      : std_logic;                     -- dma_LCD:write_write_n -> dma_lcd_write_master_write:in
	signal dma_lcd_write_master_writedata                                  : std_logic_vector(15 downto 0); -- dma_LCD:write_writedata -> mm_interconnect_0:dma_LCD_write_master_writedata
	signal mm_interconnect_0_sdram_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                             : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                          : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                              : std_logic_vector(21 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                 : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                        : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_ili9341spi_a_slave_chipselect                 : std_logic;                     -- mm_interconnect_0:ILI9341SPI_a_slave_chipselect -> ILI9341SPI:sel
	signal mm_interconnect_0_ili9341spi_a_slave_waitrequest                : std_logic;                     -- ILI9341SPI:waitreq -> mm_interconnect_0:ILI9341SPI_a_slave_waitrequest
	signal mm_interconnect_0_ili9341spi_a_slave_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ILI9341SPI_a_slave_address -> ILI9341SPI:address
	signal mm_interconnect_0_ili9341spi_a_slave_byteenable                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ILI9341SPI_a_slave_byteenable -> ILI9341SPI:ben
	signal mm_interconnect_0_ili9341spi_a_slave_write                      : std_logic;                     -- mm_interconnect_0:ILI9341SPI_a_slave_write -> ILI9341SPI:wr
	signal mm_interconnect_0_ili9341spi_a_slave_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:ILI9341SPI_a_slave_writedata -> ILI9341SPI:wrdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect        : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata          : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest       : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address           : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read              : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write             : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_ft245_avalon_slave_chipselect                 : std_logic;                     -- mm_interconnect_0:ft245_avalon_slave_chipselect -> ft245:sel
	signal mm_interconnect_0_ft245_avalon_slave_readdata                   : std_logic_vector(31 downto 0); -- ft245:rddata -> mm_interconnect_0:ft245_avalon_slave_readdata
	signal mm_interconnect_0_ft245_avalon_slave_waitrequest                : std_logic;                     -- ft245:waitreq -> mm_interconnect_0:ft245_avalon_slave_waitrequest
	signal mm_interconnect_0_ft245_avalon_slave_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:ft245_avalon_slave_address -> ft245:address
	signal mm_interconnect_0_ft245_avalon_slave_read                       : std_logic;                     -- mm_interconnect_0:ft245_avalon_slave_read -> ft245:rd
	signal mm_interconnect_0_ft245_avalon_slave_byteenable                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ft245_avalon_slave_byteenable -> ft245:ben
	signal mm_interconnect_0_ft245_avalon_slave_write                      : std_logic;                     -- mm_interconnect_0:ft245_avalon_slave_write -> ft245:wr
	signal mm_interconnect_0_ft245_avalon_slave_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:ft245_avalon_slave_writedata -> ft245:wrdata
	signal mm_interconnect_0_dma_control_port_slave_chipselect             : std_logic;                     -- mm_interconnect_0:dma_control_port_slave_chipselect -> dma:dma_ctl_chipselect
	signal mm_interconnect_0_dma_control_port_slave_readdata               : std_logic_vector(23 downto 0); -- dma:dma_ctl_readdata -> mm_interconnect_0:dma_control_port_slave_readdata
	signal mm_interconnect_0_dma_control_port_slave_address                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:dma_control_port_slave_address -> dma:dma_ctl_address
	signal mm_interconnect_0_dma_control_port_slave_write                  : std_logic;                     -- mm_interconnect_0:dma_control_port_slave_write -> mm_interconnect_0_dma_control_port_slave_write:in
	signal mm_interconnect_0_dma_control_port_slave_writedata              : std_logic_vector(23 downto 0); -- mm_interconnect_0:dma_control_port_slave_writedata -> dma:dma_ctl_writedata
	signal mm_interconnect_0_dma_lcd_control_port_slave_chipselect         : std_logic;                     -- mm_interconnect_0:dma_LCD_control_port_slave_chipselect -> dma_LCD:dma_ctl_chipselect
	signal mm_interconnect_0_dma_lcd_control_port_slave_readdata           : std_logic_vector(23 downto 0); -- dma_LCD:dma_ctl_readdata -> mm_interconnect_0:dma_LCD_control_port_slave_readdata
	signal mm_interconnect_0_dma_lcd_control_port_slave_address            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:dma_LCD_control_port_slave_address -> dma_LCD:dma_ctl_address
	signal mm_interconnect_0_dma_lcd_control_port_slave_write              : std_logic;                     -- mm_interconnect_0:dma_LCD_control_port_slave_write -> mm_interconnect_0_dma_lcd_control_port_slave_write:in
	signal mm_interconnect_0_dma_lcd_control_port_slave_writedata          : std_logic_vector(23 downto 0); -- mm_interconnect_0:dma_LCD_control_port_slave_writedata -> dma_LCD:dma_ctl_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                  : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                   : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_onchip_flash_data_readdata                    : std_logic_vector(31 downto 0); -- onchip_flash:avmm_data_readdata -> mm_interconnect_0:onchip_flash_data_readdata
	signal mm_interconnect_0_onchip_flash_data_waitrequest                 : std_logic;                     -- onchip_flash:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_data_waitrequest
	signal mm_interconnect_0_onchip_flash_data_address                     : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_flash_data_address -> onchip_flash:avmm_data_addr
	signal mm_interconnect_0_onchip_flash_data_read                        : std_logic;                     -- mm_interconnect_0:onchip_flash_data_read -> onchip_flash:avmm_data_read
	signal mm_interconnect_0_onchip_flash_data_readdatavalid               : std_logic;                     -- onchip_flash:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_data_readdatavalid
	signal mm_interconnect_0_onchip_flash_data_write                       : std_logic;                     -- mm_interconnect_0:onchip_flash_data_write -> onchip_flash:avmm_data_write
	signal mm_interconnect_0_onchip_flash_data_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_flash_data_writedata -> onchip_flash:avmm_data_writedata
	signal mm_interconnect_0_onchip_flash_data_burstcount                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_flash_data_burstcount -> onchip_flash:avmm_data_burstcount
	signal mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata           : std_logic_vector(31 downto 0); -- nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest        : std_logic;                     -- nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess        : std_logic;                     -- mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_debug_mem_slave_address            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_debug_mem_slave_read               : std_logic;                     -- mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_debug_mem_slave_write              : std_logic;                     -- mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	signal mm_interconnect_0_serialflash_epcs_control_port_chipselect      : std_logic;                     -- mm_interconnect_0:serialflash_epcs_control_port_chipselect -> serialflash:chipselect
	signal mm_interconnect_0_serialflash_epcs_control_port_readdata        : std_logic_vector(31 downto 0); -- serialflash:readdata -> mm_interconnect_0:serialflash_epcs_control_port_readdata
	signal mm_interconnect_0_serialflash_epcs_control_port_address         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:serialflash_epcs_control_port_address -> serialflash:address
	signal mm_interconnect_0_serialflash_epcs_control_port_read            : std_logic;                     -- mm_interconnect_0:serialflash_epcs_control_port_read -> mm_interconnect_0_serialflash_epcs_control_port_read:in
	signal mm_interconnect_0_serialflash_epcs_control_port_write           : std_logic;                     -- mm_interconnect_0:serialflash_epcs_control_port_write -> mm_interconnect_0_serialflash_epcs_control_port_write:in
	signal mm_interconnect_0_serialflash_epcs_control_port_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:serialflash_epcs_control_port_writedata -> serialflash:writedata
	signal mm_interconnect_0_sys_clk_timer_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_0_sys_clk_timer_s1_readdata                     : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	signal mm_interconnect_0_sys_clk_timer_s1_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_0_sys_clk_timer_s1_write                        : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_write -> mm_interconnect_0_sys_clk_timer_s1_write:in
	signal mm_interconnect_0_sys_clk_timer_s1_writedata                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_0_button_s1_readdata                            : std_logic_vector(31 downto 0); -- button:readdata -> mm_interconnect_0:button_s1_readdata
	signal mm_interconnect_0_button_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button_s1_address -> button:address
	signal mm_interconnect_0_debport_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:DEBport_s1_chipselect -> DEBport:chipselect
	signal mm_interconnect_0_debport_s1_readdata                           : std_logic_vector(31 downto 0); -- DEBport:readdata -> mm_interconnect_0:DEBport_s1_readdata
	signal mm_interconnect_0_debport_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:DEBport_s1_address -> DEBport:address
	signal mm_interconnect_0_debport_s1_write                              : std_logic;                     -- mm_interconnect_0:DEBport_s1_write -> mm_interconnect_0_debport_s1_write:in
	signal mm_interconnect_0_debport_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:DEBport_s1_writedata -> DEBport:writedata
	signal mm_interconnect_0_led_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:LED_s1_chipselect -> LED:chipselect
	signal mm_interconnect_0_led_s1_readdata                               : std_logic_vector(31 downto 0); -- LED:readdata -> mm_interconnect_0:LED_s1_readdata
	signal mm_interconnect_0_led_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LED_s1_address -> LED:address
	signal mm_interconnect_0_led_s1_write                                  : std_logic;                     -- mm_interconnect_0:LED_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:LED_s1_writedata -> LED:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- sys_clk_timer:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- serialflash:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- dma:dma_ctl_irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                        : std_logic;                     -- ft245:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                        : std_logic;                     -- dma_LCD:dma_ctl_irq -> irq_mapper:receiver5_irq
	signal nios2_gen2_irq_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2:reset_req, rst_translator:reset_req_in, serialflash:reset_req]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                              : std_logic;                     -- rst_controller_002:reset_out -> pll:reset
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal nios2_gen2_debug_reset_request_reset_ports_inv                  : std_logic;                     -- nios2_gen2_debug_reset_request_reset:inv -> [DEBport:reset_n, ILI9341SPI:reset_n, LED:reset_n, dma:system_reset_n, dma_LCD:system_reset_n, ft245:reset_n]
	signal dma_read_master_read_ports_inv                                  : std_logic;                     -- dma_read_master_read:inv -> mm_interconnect_0:dma_read_master_read
	signal dma_lcd_read_master_read_ports_inv                              : std_logic;                     -- dma_lcd_read_master_read:inv -> mm_interconnect_0:dma_LCD_read_master_read
	signal dma_write_master_write_ports_inv                                : std_logic;                     -- dma_write_master_write:inv -> mm_interconnect_0:dma_write_master_write
	signal dma_lcd_write_master_write_ports_inv                            : std_logic;                     -- dma_lcd_write_master_write:inv -> mm_interconnect_0:dma_LCD_write_master_write
	signal mm_interconnect_0_sdram_s1_read_ports_inv                       : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv    : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv   : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_dma_control_port_slave_write_ports_inv        : std_logic;                     -- mm_interconnect_0_dma_control_port_slave_write:inv -> dma:dma_ctl_write_n
	signal mm_interconnect_0_dma_lcd_control_port_slave_write_ports_inv    : std_logic;                     -- mm_interconnect_0_dma_lcd_control_port_slave_write:inv -> dma_LCD:dma_ctl_write_n
	signal mm_interconnect_0_serialflash_epcs_control_port_read_ports_inv  : std_logic;                     -- mm_interconnect_0_serialflash_epcs_control_port_read:inv -> serialflash:read_n
	signal mm_interconnect_0_serialflash_epcs_control_port_write_ports_inv : std_logic;                     -- mm_interconnect_0_serialflash_epcs_control_port_write:inv -> serialflash:write_n
	signal mm_interconnect_0_sys_clk_timer_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal mm_interconnect_0_debport_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_debport_s1_write:inv -> DEBport:write_n
	signal mm_interconnect_0_led_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> LED:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [button:reset_n, nios2_gen2:reset_n, onchip_flash:reset_n, sdram:reset_n, serialflash:reset_n, sys_clk_timer:reset_n, sysid:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> jtag_uart:rst_n

begin

	debport : component nios_DEBport
		port map (
			clk        => pll_c0_clk,                                     --                 clk.clk
			reset_n    => nios2_gen2_debug_reset_request_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_debport_s1_address,           --                  s1.address
			write_n    => mm_interconnect_0_debport_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_0_debport_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_0_debport_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_0_debport_s1_readdata,          --                    .readdata
			out_port   => deb_export                                      -- external_connection.export
		);

	ili9341spi : component ili9341_spi16
		port map (
			clk     => pll_c0_clk,                                       --       clock.clk
			reset_n => nios2_gen2_debug_reset_request_reset_ports_inv,   --       reset.reset_n
			address => mm_interconnect_0_ili9341spi_a_slave_address,     --     a_slave.address
			ben     => mm_interconnect_0_ili9341spi_a_slave_byteenable,  --            .byteenable
			sel     => mm_interconnect_0_ili9341spi_a_slave_chipselect,  --            .chipselect
			wr      => mm_interconnect_0_ili9341spi_a_slave_write,       --            .write
			wrdata  => mm_interconnect_0_ili9341spi_a_slave_writedata,   --            .writedata
			waitreq => mm_interconnect_0_ili9341spi_a_slave_waitrequest, --            .waitrequest
			cs      => lcd_cs,                                           -- conduit_end.cs
			dc      => lcd_dc,                                           --            .dc
			rstn    => lcd_rstn,                                         --            .rstn
			sclk    => lcd_sclk,                                         --            .sclk
			sdata   => lcd_sdata                                         --            .sdata
		);

	led : component nios_DEBport
		port map (
			clk        => pll_c0_clk,                                     --                 clk.clk
			reset_n    => nios2_gen2_debug_reset_request_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,               --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv,       --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,             --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,            --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,              --                    .readdata
			out_port   => led_export                                      -- external_connection.export
		);

	button : component nios_button
		port map (
			clk      => pll_c0_clk,                               --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_button_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_button_s1_readdata,     --                    .readdata
			in_port  => button_export                             -- external_connection.export
		);

	dma : component nios_dma
		port map (
			clk                => pll_c0_clk,                                               --                clk.clk
			system_reset_n     => nios2_gen2_debug_reset_request_reset_ports_inv,           --              reset.reset_n
			dma_ctl_address    => mm_interconnect_0_dma_control_port_slave_address,         -- control_port_slave.address
			dma_ctl_chipselect => mm_interconnect_0_dma_control_port_slave_chipselect,      --                   .chipselect
			dma_ctl_readdata   => mm_interconnect_0_dma_control_port_slave_readdata,        --                   .readdata
			dma_ctl_write_n    => mm_interconnect_0_dma_control_port_slave_write_ports_inv, --                   .write_n
			dma_ctl_writedata  => mm_interconnect_0_dma_control_port_slave_writedata,       --                   .writedata
			dma_ctl_irq        => irq_mapper_receiver3_irq,                                 --                irq.irq
			read_address       => dma_read_master_address,                                  --        read_master.address
			read_chipselect    => dma_read_master_chipselect,                               --                   .chipselect
			read_read_n        => dma_read_master_read,                                     --                   .read_n
			read_readdata      => dma_read_master_readdata,                                 --                   .readdata
			read_readdatavalid => dma_read_master_readdatavalid,                            --                   .readdatavalid
			read_waitrequest   => dma_read_master_waitrequest,                              --                   .waitrequest
			write_address      => dma_write_master_address,                                 --       write_master.address
			write_chipselect   => dma_write_master_chipselect,                              --                   .chipselect
			write_waitrequest  => dma_write_master_waitrequest,                             --                   .waitrequest
			write_write_n      => dma_write_master_write,                                   --                   .write_n
			write_writedata    => dma_write_master_writedata,                               --                   .writedata
			write_byteenable   => dma_write_master_byteenable                               --                   .byteenable
		);

	dma_lcd : component nios_dma_LCD
		port map (
			clk                => pll_c0_clk,                                                   --                clk.clk
			system_reset_n     => nios2_gen2_debug_reset_request_reset_ports_inv,               --              reset.reset_n
			dma_ctl_address    => mm_interconnect_0_dma_lcd_control_port_slave_address,         -- control_port_slave.address
			dma_ctl_chipselect => mm_interconnect_0_dma_lcd_control_port_slave_chipselect,      --                   .chipselect
			dma_ctl_readdata   => mm_interconnect_0_dma_lcd_control_port_slave_readdata,        --                   .readdata
			dma_ctl_write_n    => mm_interconnect_0_dma_lcd_control_port_slave_write_ports_inv, --                   .write_n
			dma_ctl_writedata  => mm_interconnect_0_dma_lcd_control_port_slave_writedata,       --                   .writedata
			dma_ctl_irq        => irq_mapper_receiver5_irq,                                     --                irq.irq
			read_address       => dma_lcd_read_master_address,                                  --        read_master.address
			read_chipselect    => dma_lcd_read_master_chipselect,                               --                   .chipselect
			read_read_n        => dma_lcd_read_master_read,                                     --                   .read_n
			read_readdata      => dma_lcd_read_master_readdata,                                 --                   .readdata
			read_readdatavalid => dma_lcd_read_master_readdatavalid,                            --                   .readdatavalid
			read_waitrequest   => dma_lcd_read_master_waitrequest,                              --                   .waitrequest
			write_address      => dma_lcd_write_master_address,                                 --       write_master.address
			write_chipselect   => dma_lcd_write_master_chipselect,                              --                   .chipselect
			write_waitrequest  => dma_lcd_write_master_waitrequest,                             --                   .waitrequest
			write_write_n      => dma_lcd_write_master_write,                                   --                   .write_n
			write_writedata    => dma_lcd_write_master_writedata,                               --                   .writedata
			write_byteenable   => dma_lcd_write_master_byteenable                               --                   .byteenable
		);

	ft245 : component ft245if2
		port map (
			address      => mm_interconnect_0_ft245_avalon_slave_address,     -- avalon_slave.address
			ben          => mm_interconnect_0_ft245_avalon_slave_byteenable,  --             .byteenable
			rd           => mm_interconnect_0_ft245_avalon_slave_read,        --             .read
			rddata       => mm_interconnect_0_ft245_avalon_slave_readdata,    --             .readdata
			sel          => mm_interconnect_0_ft245_avalon_slave_chipselect,  --             .chipselect
			waitreq      => mm_interconnect_0_ft245_avalon_slave_waitrequest, --             .waitrequest
			wr           => mm_interconnect_0_ft245_avalon_slave_write,       --             .write
			wrdata       => mm_interconnect_0_ft245_avalon_slave_writedata,   --             .writedata
			clk          => pll_c0_clk,                                       --        clock.clk
			ft_rdn       => ftdi_rdn,                                         --       export.rdn
			ft_resetn    => ftdi_resetn,                                      --             .resetn
			ft_rxdata    => ftdi_rxdata,                                      --             .rxdata
			ft_rxfn      => ftdi_rxfn,                                        --             .rxfn
			ft_txdata    => ftdi_txdata,                                      --             .txdata
			ft_txdata_oe => ftdi_txdata_oe,                                   --             .txdata_oe
			ft_txen      => ftdi_txen,                                        --             .txen
			ft_wr        => ftdi_wr,                                          --             .wr
			irq          => irq_mapper_receiver4_irq,                         --          irq.irq
			reset_n      => nios2_gen2_debug_reset_request_reset_ports_inv    --        reset.reset_n
		);

	jtag_uart : component nios_jtag_uart
		port map (
			clk            => pll_c0_clk,                                                    --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	nios2_gen2 : component nios_nios2_gen2
		port map (
			clk                                 => pll_c0_clk,                                               --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                 --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                       --                          .reset_req
			d_address                           => nios2_gen2_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                      -- custom_instruction_master.readra
		);

	onchip_flash : component altera_onchip_flash
		generic map (
			INIT_FILENAME                       => "",
			INIT_FILENAME_SIM                   => "",
			DEVICE_FAMILY                       => "MAX 10",
			PART_NAME                           => "10M08DAF484C8GES",
			DEVICE_ID                           => "08",
			SECTOR1_START_ADDR                  => 0,
			SECTOR1_END_ADDR                    => 4095,
			SECTOR2_START_ADDR                  => 4096,
			SECTOR2_END_ADDR                    => 8191,
			SECTOR3_START_ADDR                  => 0,
			SECTOR3_END_ADDR                    => 0,
			SECTOR4_START_ADDR                  => 0,
			SECTOR4_END_ADDR                    => 0,
			SECTOR5_START_ADDR                  => 0,
			SECTOR5_END_ADDR                    => 0,
			MIN_VALID_ADDR                      => 0,
			MAX_VALID_ADDR                      => 8191,
			MIN_UFM_VALID_ADDR                  => 0,
			MAX_UFM_VALID_ADDR                  => 8191,
			SECTOR1_MAP                         => 1,
			SECTOR2_MAP                         => 2,
			SECTOR3_MAP                         => 0,
			SECTOR4_MAP                         => 0,
			SECTOR5_MAP                         => 0,
			ADDR_RANGE1_END_ADDR                => 8191,
			ADDR_RANGE2_END_ADDR                => 8191,
			ADDR_RANGE1_OFFSET                  => 512,
			ADDR_RANGE2_OFFSET                  => 0,
			ADDR_RANGE3_OFFSET                  => 0,
			AVMM_DATA_ADDR_WIDTH                => 13,
			AVMM_DATA_DATA_WIDTH                => 32,
			AVMM_DATA_BURSTCOUNT_WIDTH          => 4,
			SECTOR_READ_PROTECTION_MODE         => 28,
			FLASH_SEQ_READ_DATA_COUNT           => 2,
			FLASH_ADDR_ALIGNMENT_BITS           => 1,
			FLASH_READ_CYCLE_MAX_INDEX          => 4,
			FLASH_RESET_CYCLE_MAX_INDEX         => 12,
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  => 60,
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX => 17500000,
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX => 15250,
			PARALLEL_MODE                       => true,
			READ_AND_WRITE_MODE                 => true,
			WRAPPING_BURST_MODE                 => false,
			IS_DUAL_BOOT                        => "False",
			IS_ERAM_SKIP                        => "False",
			IS_COMPRESSED_IMAGE                 => "False"
		)
		port map (
			clock                   => pll_c0_clk,                                        --    clk.clk
			reset_n                 => rst_controller_reset_out_reset_ports_inv,          -- nreset.reset_n
			avmm_data_addr          => mm_interconnect_0_onchip_flash_data_address,       --   data.address
			avmm_data_read          => mm_interconnect_0_onchip_flash_data_read,          --       .read
			avmm_data_writedata     => mm_interconnect_0_onchip_flash_data_writedata,     --       .writedata
			avmm_data_write         => mm_interconnect_0_onchip_flash_data_write,         --       .write
			avmm_data_readdata      => mm_interconnect_0_onchip_flash_data_readdata,      --       .readdata
			avmm_data_waitrequest   => mm_interconnect_0_onchip_flash_data_waitrequest,   --       .waitrequest
			avmm_data_readdatavalid => mm_interconnect_0_onchip_flash_data_readdatavalid, --       .readdatavalid
			avmm_data_burstcount    => mm_interconnect_0_onchip_flash_data_burstcount,    --       .burstcount
			avmm_csr_addr           => open,                                              --    csr.address
			avmm_csr_read           => open,                                              --       .read
			avmm_csr_writedata      => open,                                              --       .writedata
			avmm_csr_write          => open,                                              --       .write
			avmm_csr_readdata       => open                                               --       .readdata
		);

	pll : component nios_pll
		port map (
			clk                => clk_clk,                            --       inclk_interface.clk
			reset              => rst_controller_002_reset_out_reset, -- inclk_interface_reset.reset
			read               => open,                               --             pll_slave.read
			write              => open,                               --                      .write
			address            => open,                               --                      .address
			readdata           => open,                               --                      .readdata
			writedata          => open,                               --                      .writedata
			c0                 => pll_c0_clk,                         --                    c0.clk
			c1                 => sd_clk,                             --                    c1.clk
			c2                 => sys_clk,                            --                    c2.clk
			c3                 => pdm_clk,                            --                    c3.clk
			c4                 => log_clk,                            --                    c4.clk
			locked             => pll_lock_export,                    --        locked_conduit.export
			scandone           => open,                               --           (terminated)
			scandataout        => open,                               --           (terminated)
			areset             => '0',                                --           (terminated)
			phasedone          => open,                               --           (terminated)
			phasecounterselect => "000",                              --           (terminated)
			phaseupdown        => '0',                                --           (terminated)
			phasestep          => '0',                                --           (terminated)
			scanclk            => '0',                                --           (terminated)
			scanclkena         => '0',                                --           (terminated)
			scandata           => '0',                                --           (terminated)
			configupdate       => '0'                                 --           (terminated)
		);

	sdram : component nios_sdram
		port map (
			clk            => pll_c0_clk,                                      --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	serialflash : component nios_serialflash
		port map (
			clk        => pll_c0_clk,                                                      --               clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			reset_req  => rst_controller_reset_out_reset_req,                              --                  .reset_req
			address    => mm_interconnect_0_serialflash_epcs_control_port_address,         -- epcs_control_port.address
			chipselect => mm_interconnect_0_serialflash_epcs_control_port_chipselect,      --                  .chipselect
			read_n     => mm_interconnect_0_serialflash_epcs_control_port_read_ports_inv,  --                  .read_n
			readdata   => mm_interconnect_0_serialflash_epcs_control_port_readdata,        --                  .readdata
			write_n    => mm_interconnect_0_serialflash_epcs_control_port_write_ports_inv, --                  .write_n
			writedata  => mm_interconnect_0_serialflash_epcs_control_port_writedata,       --                  .writedata
			irq        => irq_mapper_receiver2_irq,                                        --               irq.irq
			dclk       => sflash_dclk,                                                     --          external.export
			sce        => sflash_sce,                                                      --                  .export
			sdo        => sflash_sdo,                                                      --                  .export
			data0      => sflash_data0                                                     --                  .export
		);

	sys_clk_timer : component nios_sys_clk_timer
		port map (
			clk        => pll_c0_clk,                                         --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           -- reset.reset_n
			address    => mm_interconnect_0_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                            --   irq.irq
		);

	sysid : component nios_sysid
		port map (
			clock    => pll_c0_clk,                                       --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component nios_mm_interconnect_0
		port map (
			pll_c0_clk                                            => pll_c0_clk,                                                 --                                          pll_c0.clk
			av_wr_master_0_reset_sink_reset_bridge_in_reset_reset => nios2_gen2_debug_reset_request_reset,                       -- av_wr_master_0_reset_sink_reset_bridge_in_reset.reset
			jtag_uart_reset_reset_bridge_in_reset_reset           => rst_controller_001_reset_out_reset,                         --           jtag_uart_reset_reset_bridge_in_reset.reset
			nios2_gen2_reset_reset_bridge_in_reset_reset          => rst_controller_reset_out_reset,                             --          nios2_gen2_reset_reset_bridge_in_reset.reset
			av_wr_master_0_avalon_master_address                  => amwr_address,                                               --                    av_wr_master_0_avalon_master.address
			av_wr_master_0_avalon_master_waitrequest              => amwr_waitrequest,                                           --                                                .waitrequest
			av_wr_master_0_avalon_master_burstcount               => amwr_burstcount,                                            --                                                .burstcount
			av_wr_master_0_avalon_master_byteenable               => amwr_byteenable,                                            --                                                .byteenable
			av_wr_master_0_avalon_master_write                    => amwr_write,                                                 --                                                .write
			av_wr_master_0_avalon_master_writedata                => amwr_writedata,                                             --                                                .writedata
			dma_read_master_address                               => dma_read_master_address,                                    --                                 dma_read_master.address
			dma_read_master_waitrequest                           => dma_read_master_waitrequest,                                --                                                .waitrequest
			dma_read_master_chipselect                            => dma_read_master_chipselect,                                 --                                                .chipselect
			dma_read_master_read                                  => dma_read_master_read_ports_inv,                             --                                                .read
			dma_read_master_readdata                              => dma_read_master_readdata,                                   --                                                .readdata
			dma_read_master_readdatavalid                         => dma_read_master_readdatavalid,                              --                                                .readdatavalid
			dma_write_master_address                              => dma_write_master_address,                                   --                                dma_write_master.address
			dma_write_master_waitrequest                          => dma_write_master_waitrequest,                               --                                                .waitrequest
			dma_write_master_byteenable                           => dma_write_master_byteenable,                                --                                                .byteenable
			dma_write_master_chipselect                           => dma_write_master_chipselect,                                --                                                .chipselect
			dma_write_master_write                                => dma_write_master_write_ports_inv,                           --                                                .write
			dma_write_master_writedata                            => dma_write_master_writedata,                                 --                                                .writedata
			dma_LCD_read_master_address                           => dma_lcd_read_master_address,                                --                             dma_LCD_read_master.address
			dma_LCD_read_master_waitrequest                       => dma_lcd_read_master_waitrequest,                            --                                                .waitrequest
			dma_LCD_read_master_chipselect                        => dma_lcd_read_master_chipselect,                             --                                                .chipselect
			dma_LCD_read_master_read                              => dma_lcd_read_master_read_ports_inv,                         --                                                .read
			dma_LCD_read_master_readdata                          => dma_lcd_read_master_readdata,                               --                                                .readdata
			dma_LCD_read_master_readdatavalid                     => dma_lcd_read_master_readdatavalid,                          --                                                .readdatavalid
			dma_LCD_write_master_address                          => dma_lcd_write_master_address,                               --                            dma_LCD_write_master.address
			dma_LCD_write_master_waitrequest                      => dma_lcd_write_master_waitrequest,                           --                                                .waitrequest
			dma_LCD_write_master_byteenable                       => dma_lcd_write_master_byteenable,                            --                                                .byteenable
			dma_LCD_write_master_chipselect                       => dma_lcd_write_master_chipselect,                            --                                                .chipselect
			dma_LCD_write_master_write                            => dma_lcd_write_master_write_ports_inv,                       --                                                .write
			dma_LCD_write_master_writedata                        => dma_lcd_write_master_writedata,                             --                                                .writedata
			nios2_gen2_data_master_address                        => nios2_gen2_data_master_address,                             --                          nios2_gen2_data_master.address
			nios2_gen2_data_master_waitrequest                    => nios2_gen2_data_master_waitrequest,                         --                                                .waitrequest
			nios2_gen2_data_master_byteenable                     => nios2_gen2_data_master_byteenable,                          --                                                .byteenable
			nios2_gen2_data_master_read                           => nios2_gen2_data_master_read,                                --                                                .read
			nios2_gen2_data_master_readdata                       => nios2_gen2_data_master_readdata,                            --                                                .readdata
			nios2_gen2_data_master_write                          => nios2_gen2_data_master_write,                               --                                                .write
			nios2_gen2_data_master_writedata                      => nios2_gen2_data_master_writedata,                           --                                                .writedata
			nios2_gen2_data_master_debugaccess                    => nios2_gen2_data_master_debugaccess,                         --                                                .debugaccess
			nios2_gen2_instruction_master_address                 => nios2_gen2_instruction_master_address,                      --                   nios2_gen2_instruction_master.address
			nios2_gen2_instruction_master_waitrequest             => nios2_gen2_instruction_master_waitrequest,                  --                                                .waitrequest
			nios2_gen2_instruction_master_read                    => nios2_gen2_instruction_master_read,                         --                                                .read
			nios2_gen2_instruction_master_readdata                => nios2_gen2_instruction_master_readdata,                     --                                                .readdata
			button_s1_address                                     => mm_interconnect_0_button_s1_address,                        --                                       button_s1.address
			button_s1_readdata                                    => mm_interconnect_0_button_s1_readdata,                       --                                                .readdata
			DEBport_s1_address                                    => mm_interconnect_0_debport_s1_address,                       --                                      DEBport_s1.address
			DEBport_s1_write                                      => mm_interconnect_0_debport_s1_write,                         --                                                .write
			DEBport_s1_readdata                                   => mm_interconnect_0_debport_s1_readdata,                      --                                                .readdata
			DEBport_s1_writedata                                  => mm_interconnect_0_debport_s1_writedata,                     --                                                .writedata
			DEBport_s1_chipselect                                 => mm_interconnect_0_debport_s1_chipselect,                    --                                                .chipselect
			dma_control_port_slave_address                        => mm_interconnect_0_dma_control_port_slave_address,           --                          dma_control_port_slave.address
			dma_control_port_slave_write                          => mm_interconnect_0_dma_control_port_slave_write,             --                                                .write
			dma_control_port_slave_readdata                       => mm_interconnect_0_dma_control_port_slave_readdata,          --                                                .readdata
			dma_control_port_slave_writedata                      => mm_interconnect_0_dma_control_port_slave_writedata,         --                                                .writedata
			dma_control_port_slave_chipselect                     => mm_interconnect_0_dma_control_port_slave_chipselect,        --                                                .chipselect
			dma_LCD_control_port_slave_address                    => mm_interconnect_0_dma_lcd_control_port_slave_address,       --                      dma_LCD_control_port_slave.address
			dma_LCD_control_port_slave_write                      => mm_interconnect_0_dma_lcd_control_port_slave_write,         --                                                .write
			dma_LCD_control_port_slave_readdata                   => mm_interconnect_0_dma_lcd_control_port_slave_readdata,      --                                                .readdata
			dma_LCD_control_port_slave_writedata                  => mm_interconnect_0_dma_lcd_control_port_slave_writedata,     --                                                .writedata
			dma_LCD_control_port_slave_chipselect                 => mm_interconnect_0_dma_lcd_control_port_slave_chipselect,    --                                                .chipselect
			ft245_avalon_slave_address                            => mm_interconnect_0_ft245_avalon_slave_address,               --                              ft245_avalon_slave.address
			ft245_avalon_slave_write                              => mm_interconnect_0_ft245_avalon_slave_write,                 --                                                .write
			ft245_avalon_slave_read                               => mm_interconnect_0_ft245_avalon_slave_read,                  --                                                .read
			ft245_avalon_slave_readdata                           => mm_interconnect_0_ft245_avalon_slave_readdata,              --                                                .readdata
			ft245_avalon_slave_writedata                          => mm_interconnect_0_ft245_avalon_slave_writedata,             --                                                .writedata
			ft245_avalon_slave_byteenable                         => mm_interconnect_0_ft245_avalon_slave_byteenable,            --                                                .byteenable
			ft245_avalon_slave_waitrequest                        => mm_interconnect_0_ft245_avalon_slave_waitrequest,           --                                                .waitrequest
			ft245_avalon_slave_chipselect                         => mm_interconnect_0_ft245_avalon_slave_chipselect,            --                                                .chipselect
			ILI9341SPI_a_slave_address                            => mm_interconnect_0_ili9341spi_a_slave_address,               --                              ILI9341SPI_a_slave.address
			ILI9341SPI_a_slave_write                              => mm_interconnect_0_ili9341spi_a_slave_write,                 --                                                .write
			ILI9341SPI_a_slave_writedata                          => mm_interconnect_0_ili9341spi_a_slave_writedata,             --                                                .writedata
			ILI9341SPI_a_slave_byteenable                         => mm_interconnect_0_ili9341spi_a_slave_byteenable,            --                                                .byteenable
			ILI9341SPI_a_slave_waitrequest                        => mm_interconnect_0_ili9341spi_a_slave_waitrequest,           --                                                .waitrequest
			ILI9341SPI_a_slave_chipselect                         => mm_interconnect_0_ili9341spi_a_slave_chipselect,            --                                                .chipselect
			jtag_uart_avalon_jtag_slave_address                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,      --                     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,        --                                                .write
			jtag_uart_avalon_jtag_slave_read                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,         --                                                .read
			jtag_uart_avalon_jtag_slave_readdata                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,     --                                                .readdata
			jtag_uart_avalon_jtag_slave_writedata                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,    --                                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,  --                                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,   --                                                .chipselect
			LED_s1_address                                        => mm_interconnect_0_led_s1_address,                           --                                          LED_s1.address
			LED_s1_write                                          => mm_interconnect_0_led_s1_write,                             --                                                .write
			LED_s1_readdata                                       => mm_interconnect_0_led_s1_readdata,                          --                                                .readdata
			LED_s1_writedata                                      => mm_interconnect_0_led_s1_writedata,                         --                                                .writedata
			LED_s1_chipselect                                     => mm_interconnect_0_led_s1_chipselect,                        --                                                .chipselect
			nios2_gen2_debug_mem_slave_address                    => mm_interconnect_0_nios2_gen2_debug_mem_slave_address,       --                      nios2_gen2_debug_mem_slave.address
			nios2_gen2_debug_mem_slave_write                      => mm_interconnect_0_nios2_gen2_debug_mem_slave_write,         --                                                .write
			nios2_gen2_debug_mem_slave_read                       => mm_interconnect_0_nios2_gen2_debug_mem_slave_read,          --                                                .read
			nios2_gen2_debug_mem_slave_readdata                   => mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata,      --                                                .readdata
			nios2_gen2_debug_mem_slave_writedata                  => mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata,     --                                                .writedata
			nios2_gen2_debug_mem_slave_byteenable                 => mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable,    --                                                .byteenable
			nios2_gen2_debug_mem_slave_waitrequest                => mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest,   --                                                .waitrequest
			nios2_gen2_debug_mem_slave_debugaccess                => mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess,   --                                                .debugaccess
			onchip_flash_data_address                             => mm_interconnect_0_onchip_flash_data_address,                --                               onchip_flash_data.address
			onchip_flash_data_write                               => mm_interconnect_0_onchip_flash_data_write,                  --                                                .write
			onchip_flash_data_read                                => mm_interconnect_0_onchip_flash_data_read,                   --                                                .read
			onchip_flash_data_readdata                            => mm_interconnect_0_onchip_flash_data_readdata,               --                                                .readdata
			onchip_flash_data_writedata                           => mm_interconnect_0_onchip_flash_data_writedata,              --                                                .writedata
			onchip_flash_data_burstcount                          => mm_interconnect_0_onchip_flash_data_burstcount,             --                                                .burstcount
			onchip_flash_data_readdatavalid                       => mm_interconnect_0_onchip_flash_data_readdatavalid,          --                                                .readdatavalid
			onchip_flash_data_waitrequest                         => mm_interconnect_0_onchip_flash_data_waitrequest,            --                                                .waitrequest
			pdm_s0_address                                        => as_pdm_address,                                             --                                          pdm_s0.address
			pdm_s0_write                                          => as_pdm_write,                                               --                                                .write
			pdm_s0_read                                           => as_pdm_read,                                                --                                                .read
			pdm_s0_readdata                                       => as_pdm_readdata,                                            --                                                .readdata
			pdm_s0_writedata                                      => as_pdm_writedata,                                           --                                                .writedata
			pdm_s0_byteenable                                     => as_pdm_byteenable,                                          --                                                .byteenable
			pdm_s0_chipselect                                     => as_pdm_chipselect,                                          --                                                .chipselect
			sdram_s1_address                                      => mm_interconnect_0_sdram_s1_address,                         --                                        sdram_s1.address
			sdram_s1_write                                        => mm_interconnect_0_sdram_s1_write,                           --                                                .write
			sdram_s1_read                                         => mm_interconnect_0_sdram_s1_read,                            --                                                .read
			sdram_s1_readdata                                     => mm_interconnect_0_sdram_s1_readdata,                        --                                                .readdata
			sdram_s1_writedata                                    => mm_interconnect_0_sdram_s1_writedata,                       --                                                .writedata
			sdram_s1_byteenable                                   => mm_interconnect_0_sdram_s1_byteenable,                      --                                                .byteenable
			sdram_s1_readdatavalid                                => mm_interconnect_0_sdram_s1_readdatavalid,                   --                                                .readdatavalid
			sdram_s1_waitrequest                                  => mm_interconnect_0_sdram_s1_waitrequest,                     --                                                .waitrequest
			sdram_s1_chipselect                                   => mm_interconnect_0_sdram_s1_chipselect,                      --                                                .chipselect
			serialflash_epcs_control_port_address                 => mm_interconnect_0_serialflash_epcs_control_port_address,    --                   serialflash_epcs_control_port.address
			serialflash_epcs_control_port_write                   => mm_interconnect_0_serialflash_epcs_control_port_write,      --                                                .write
			serialflash_epcs_control_port_read                    => mm_interconnect_0_serialflash_epcs_control_port_read,       --                                                .read
			serialflash_epcs_control_port_readdata                => mm_interconnect_0_serialflash_epcs_control_port_readdata,   --                                                .readdata
			serialflash_epcs_control_port_writedata               => mm_interconnect_0_serialflash_epcs_control_port_writedata,  --                                                .writedata
			serialflash_epcs_control_port_chipselect              => mm_interconnect_0_serialflash_epcs_control_port_chipselect, --                                                .chipselect
			sys_clk_timer_s1_address                              => mm_interconnect_0_sys_clk_timer_s1_address,                 --                                sys_clk_timer_s1.address
			sys_clk_timer_s1_write                                => mm_interconnect_0_sys_clk_timer_s1_write,                   --                                                .write
			sys_clk_timer_s1_readdata                             => mm_interconnect_0_sys_clk_timer_s1_readdata,                --                                                .readdata
			sys_clk_timer_s1_writedata                            => mm_interconnect_0_sys_clk_timer_s1_writedata,               --                                                .writedata
			sys_clk_timer_s1_chipselect                           => mm_interconnect_0_sys_clk_timer_s1_chipselect,              --                                                .chipselect
			sysid_control_slave_address                           => mm_interconnect_0_sysid_control_slave_address,              --                             sysid_control_slave.address
			sysid_control_slave_readdata                          => mm_interconnect_0_sysid_control_slave_readdata              --                                                .readdata
		);

	irq_mapper : component nios_irq_mapper
		port map (
			clk           => pll_c0_clk,                     --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,       -- receiver5.irq
			sender_irq    => nios2_gen2_irq_irq              --    sender.irq
		);

	rst_controller : component nios_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,              -- reset_in0.reset
			reset_in1      => nios2_gen2_debug_reset_request_reset, -- reset_in1.reset
			clk            => pll_c0_clk,                           --       clk.clk
			reset_out      => rst_controller_reset_out_reset,       -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,   --          .reset_req
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_001 : component nios_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_c0_clk,                         --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component nios_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	nios2_gen2_debug_reset_request_reset_ports_inv <= not nios2_gen2_debug_reset_request_reset;

	dma_read_master_read_ports_inv <= not dma_read_master_read;

	dma_lcd_read_master_read_ports_inv <= not dma_lcd_read_master_read;

	dma_write_master_write_ports_inv <= not dma_write_master_write;

	dma_lcd_write_master_write_ports_inv <= not dma_lcd_write_master_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_dma_control_port_slave_write_ports_inv <= not mm_interconnect_0_dma_control_port_slave_write;

	mm_interconnect_0_dma_lcd_control_port_slave_write_ports_inv <= not mm_interconnect_0_dma_lcd_control_port_slave_write;

	mm_interconnect_0_serialflash_epcs_control_port_read_ports_inv <= not mm_interconnect_0_serialflash_epcs_control_port_read;

	mm_interconnect_0_serialflash_epcs_control_port_write_ports_inv <= not mm_interconnect_0_serialflash_epcs_control_port_write;

	mm_interconnect_0_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_clk_timer_s1_write;

	mm_interconnect_0_debport_s1_write_ports_inv <= not mm_interconnect_0_debport_s1_write;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of nios
